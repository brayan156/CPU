module Character_manager(input logic clk,reset,
								input logic[7:0] char_data[255:0],
								input logic[7:0] char_data_coded[255:0],
								output logic [7:0] data[703:0]);

								
	logic fin;							
								
	always_ff @(posedge clk, posedge reset) begin
		if (reset) fin=0;
		else begin
		
		
		
		end
		
	end
								
								
	assign data[63:0]='{8'h54,8'h65,8'h78,8'h74,8'h6f,8'h20,8'h63,8'h6f,8'h64,8'h69,8'h66,8'h69,8'h63,8'h61,8'h64,8'h6f,8'h3a,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20};
	assign data[319:64]=char_data_coded;
	assign data[383:320]='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20};
	assign data[447:384]={8'h54,8'h65,8'h78,8'h74,8'h6f,8'h20,8'h64,8'h65,8'h63,8'h6f,8'h64,8'h69,8'h66,8'h69,8'h63,8'h61,8'h64,8'h6f,8'h20,8'h63,8'h6f,8'h6e,8'h3a,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20};
	assign data[703:448]=char_data;
	
endmodule 