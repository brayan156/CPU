module Character_manager(input logic clk,reset,swxor2,swxor1,swxor0,swxor,swnot,swadd,swinit,
								input logic[7:0] char_data[255:0],
								input logic[7:0] char_data_coded[255:0],
								output logic [7:0] data[703:0]);

								
	logic fin;							
	logic [7:0] decoded_line[63:0];					
	always_ff @(posedge clk, posedge reset) begin
		if (reset) begin fin=0;
			decoded_line='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54};	
		end
		else begin
			if (swinit) begin fin=1; end;
			if (fin) data[703:448]= char_data; else data[703:448]='{256{8'h20}};
			if (!fin)begin
				if (swxor)
					case ({swxor2,swxor1,swxor0})
					3'b000 : decoded_line ='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h30,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b001 : decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h31,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b010 : decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h32,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b011 : decoded_line ='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h33,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b100 : decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h34,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b101 : decoded_line ='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h35,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b110 : decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h36,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					3'b111 : decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h37,8'h20,8'h52,8'h4f,8'h58,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54
};
					endcase
				else if (swnot) decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h54,8'h4f,8'h4e,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54};
				else if (swadd) decoded_line = '{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h44,8'h44,8'h41,8'h20,8'h6f,8'h64,8'h6f,8'h74,8'h65,8'h6d,8'h20,8'h6e,8'h6f,8'h63,8'h20,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54};
				else decoded_line='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h65,8'h64,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54};	
		
				end	
		end
		
	end
								
								
	assign data[63:0]='{8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h20,8'h3a,8'h6f,8'h64,8'h61,8'h63,8'h69,8'h66,8'h69,8'h64,8'h6f,8'h63,8'h20,8'h6f,8'h74,8'h78,8'h65,8'h54};
	assign data[319:64]=char_data_coded;
	assign data[383:320]='{64{8'h20}};
	assign data[447:384]= decoded_line;

	
endmodule 